`ifndef __TOP_DEFINE_VH
`define __TOP_DEFINE_VH 1

`define WIDTH_DEF 32
`define DEPTH_DEF 16

`endif